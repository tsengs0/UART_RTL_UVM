//`include "uart_config.sv"
`include "uartTX_seq_item.sv"
`include "sequence/reset_clk_seq.sv"
`include "sequence/variable_baud_seq.sv"
`include "uartTX_driver.sv"
`include "uartTX_monitor.sv"
`include "uartTX_agent.sv"
`include "uart_scoreboard.sv"
`include "uart_env.sv"
`include "uart_test.sv"