typedef enum bit [1:0] {
    reset_active = 0,
    random_baud = 1
} operation_mode;